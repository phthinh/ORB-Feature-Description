module Atan2_Decoder(in, index1, index2);

parameter WIDTH = 16;
parameter WIDTH_INDEX = 5;

input [WIDTH-1:0] in;
output reg [WIDTH_INDEX-1:0] index1;
output wire [WIDTH_INDEX-1:0] index2;

always @* begin
    case(in)
	25'b1_1111_1111_1111_1111_1111_1111: index1 = 5'b00000;
	25'b1_1111_1111_1111_1111_1111_1110: index1 = 5'b00000;
	25'b1_1111_1111_1111_1111_1111_1100: index1 = 5'b00001;
	25'b1_1111_1111_1111_1111_1111_1000: index1 = 5'b00010;
	25'b1_1111_1111_1111_1111_1111_0000: index1 = 5'b00011;
	25'b1_1111_1111_1111_1111_1110_0000: index1 = 5'b00100;
	25'b1_1111_1111_1111_1111_1100_0000: index1 = 5'b00101;
	25'b1_1111_1111_1111_1111_1000_0000: index1 = 5'b00110;
	25'b1_1111_1111_1111_1111_0000_0000: index1 = 5'b00111;
	25'b1_1111_1111_1111_1110_0000_0000: index1 = 5'b01000;
	25'b1_1111_1111_1111_1100_0000_0000: index1 = 5'b01001;
	25'b1_1111_1111_1111_1000_0000_0000: index1 = 5'b01010;
	25'b1_1111_1111_1111_0000_0000_0000: index1 = 5'b01011;
	25'b1_1111_1111_1110_0000_0000_0000: index1 = 5'b01100;
	25'b1_1111_1111_1100_0000_0000_0000: index1 = 5'b01101;
	25'b1_1111_1111_1000_0000_0000_0000: index1 = 5'b01110;
	25'b1_1111_1111_0000_0000_0000_0000: index1 = 5'b01111;
	25'b1_1111_1110_0000_0000_0000_0000: index1 = 5'b10000;
	25'b1_1111_1100_0000_0000_0000_0000: index1 = 5'b10001;
	25'b1_1111_1000_0000_0000_0000_0000: index1 = 5'b10010;
	25'b1_1111_0000_0000_0000_0000_0000: index1 = 5'b10011;
	25'b1_1110_0000_0000_0000_0000_0000: index1 = 5'b10100;
	25'b1_1100_0000_0000_0000_0000_0000: index1 = 5'b10101;
	25'b1_1000_0000_0000_0000_0000_0000: index1 = 5'b10110;
	25'b1_0000_0000_0000_0000_0000_0000: index1 = 5'b10111;
	25'b0_0000_0000_0000_0000_0000_0000: index1 = 5'b11000;
	default: index1 = 5'bxxxxx;
    endcase
end

assign index2 = (|in == 1'b0) || (&in == 1'b1) ? index1: index1 + 1;

//always @* begin
//    case(in)
//	25'b1_1111_1111_1111_1111_1111_1111: index2 = 5'b00000;
//	25'b1_1111_1111_1111_1111_1111_1110: index2 = 5'b00001;
//	25'b1_1111_1111_1111_1111_1111_1100: index2 = 5'b00010;
//	25'b1_1111_1111_1111_1111_1111_1000: index2 = 5'b00011;
//	25'b1_1111_1111_1111_1111_1111_0000: index2 = 5'b00100;
//	25'b1_1111_1111_1111_1111_1110_0000: index2 = 5'b00101;
//	25'b1_1111_1111_1111_1111_1100_0000: index2 = 5'b00110;
//	25'b1_1111_1111_1111_1111_1000_0000: index2 = 5'b00111;
//	25'b1_1111_1111_1111_1111_0000_0000: index2 = 5'b01000;
//	25'b1_1111_1111_1111_1110_0000_0000: index2 = 5'b01001;
//	25'b1_1111_1111_1111_1100_0000_0000: index2 = 5'b01010;
//	25'b1_1111_1111_1111_1000_0000_0000: index2 = 5'b01011;
//	25'b1_1111_1111_1111_0000_0000_0000: index2 = 5'b01100;
//	25'b1_1111_1111_1110_0000_0000_0000: index2 = 5'b01101;
//	25'b1_1111_1111_1100_0000_0000_0000: index2 = 5'b01110;
//	25'b1_1111_1111_1000_0000_0000_0000: index2 = 5'b01111;
//	25'b1_1111_1111_0000_0000_0000_0000: index2 = 5'b10000;
//	25'b1_1111_1110_0000_0000_0000_0000: index2 = 5'b10001;
//	25'b1_1111_1100_0000_0000_0000_0000: index2 = 5'b10010;
//	25'b1_1111_1000_0000_0000_0000_0000: index2 = 5'b10011;
//	25'b1_1111_0000_0000_0000_0000_0000: index2 = 5'b10100;
//	25'b1_1110_0000_0000_0000_0000_0000: index2 = 5'b10101;
//	25'b1_1100_0000_0000_0000_0000_0000: index2 = 5'b10110;
//	25'b1_1000_0000_0000_0000_0000_0000: index2 = 5'b10111;
//	25'b1_0000_0000_0000_0000_0000_0000: index2 = 5'b11000;
//	25'b0_0000_0000_0000_0000_0000_0000: index2 = 5'b11000;
//	default: index2 = 5'bxxxxx;
//    endcase
//end
//

endmodule