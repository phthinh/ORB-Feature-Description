module MultY_connect(in0,  in1,  in2,  in3,  in4,  in5,  in6,  in7,  in8, in9, 
							in10, in11, in12, in13, in14, in15, in16, in17, in18, 
							out); 
 
parameter BW_XCOS = 16;

input signed [BW_XCOS-1:0] in0; 
input signed [BW_XCOS-1:0] in1; 
input signed [BW_XCOS-1:0] in2;  
input signed [BW_XCOS-1:0] in3;  
input signed [BW_XCOS-1:0] in4;  
input signed [BW_XCOS-1:0] in5;  
input signed [BW_XCOS-1:0] in6;  
input signed [BW_XCOS-1:0] in7;  
input signed [BW_XCOS-1:0] in8;  
input signed [BW_XCOS-1:0] in9;  
input signed [BW_XCOS-1:0] in10;  
input signed [BW_XCOS-1:0] in11;  
input signed [BW_XCOS-1:0] in12;  
input signed [BW_XCOS-1:0] in13;  
input signed [BW_XCOS-1:0] in14;  
input signed [BW_XCOS-1:0] in15;  
input signed [BW_XCOS-1:0] in16;
input signed [BW_XCOS-1:0] in17;
input signed [BW_XCOS-1:0] in18;

output [512*BW_XCOS-1:0] out; 

wire signed [BW_XCOS-1:0] res [0:511]; 

wire signed [BW_XCOS-1:0] neg0, neg1, neg2, neg3, neg4, neg5,neg6, neg7, neg8, neg9, neg10, 
	neg11, neg12, neg13, neg14, neg15, neg16, neg17, neg18; 

assign neg0=-in0;
assign neg1=-in1; 
assign neg2=-in2; 
assign neg3=-in3; 
assign neg4=-in4; 
assign neg5=-in5; 
assign neg6=-in6; 
assign neg7=-in7; 
assign neg8=-in8; 
assign neg9=-in9; 
assign neg10=-in10; 
assign neg11=-in11; 
assign neg12=-in12; 
assign neg13=-in13; 
assign neg14=-in14; 
assign neg15=-in15; 
assign neg16=-in16;
assign neg17=-in17;
assign neg18=-in18;

//Generating to assign 512 outputs of multiplication == 
assign res[0]=neg3; 
assign res[1]=in5; 
assign res[2]=in2; 
assign res[3]=neg12; 
assign res[4]=in9; 
assign res[5]=in2; 
assign res[6]=neg12; 
assign res[7]=neg13; 
assign res[8]=neg13; 
assign res[9]=in12; 
assign res[10]=neg7; 
assign res[11]=in6; 
assign res[12]=neg10; 
assign res[13]=neg4; 
assign res[14]=neg13; 
assign res[15]=neg8; 
assign res[16]=neg3; 
assign res[17]=neg9; 
assign res[18]=in4; 
assign res[19]=in9; 
assign res[20]=neg8; 
assign res[21]=neg9; 
assign res[22]=in7; 
assign res[23]=in12; 
assign res[24]=in7; 
assign res[25]=in6; 
assign res[26]=neg5; 
assign res[27]=neg0; 
assign res[28]=in2; 
assign res[29]=neg3; 
assign res[30]=neg0; 
assign res[31]=in5; 
assign res[32]=neg6; 
assign res[33]=neg1; 
assign res[34]=in6; 
assign res[35]=in12; 
assign res[36]=neg13; 
assign res[37]=neg8; 
assign res[38]=neg13; 
assign res[39]=neg8; 
assign res[40]=in7; 
assign res[41]=in1; 
assign res[42]=neg3; 
assign res[43]=neg3; 
assign res[44]=neg7; 
assign res[45]=in12; 
assign res[46]=neg7; 
assign res[47]=neg2; 
assign res[48]=in11; 
assign res[49]=neg10; 
assign res[50]=in12; 
assign res[51]=in10; 
assign res[52]=in3; 
assign res[53]=neg3; 
assign res[54]=in2; 
assign res[55]=in7; 
assign res[56]=neg12; 
assign res[57]=in11; 
assign res[58]=neg12; 
assign res[59]=neg7; 
assign res[60]=neg6; 
assign res[61]=neg1; 
assign res[62]=neg0; 
assign res[63]=neg5; 
assign res[64]=in11; 
assign res[65]=neg13; 
assign res[66]=in7; 
assign res[67]=in12; 
assign res[68]=neg1; 
assign res[69]=in4; 
assign res[70]=neg12; 
assign res[71]=in7; 
assign res[72]=neg5; 
assign res[73]=neg10; 
assign res[74]=in11; 
assign res[75]=in12; 
assign res[76]=neg8; 
assign res[77]=neg13; 
assign res[78]=neg2; 
assign res[79]=in2; 
assign res[80]=neg2; 
assign res[81]=in3; 
assign res[82]=in9; 
assign res[83]=neg9; 
assign res[84]=in12; 
assign res[85]=in7; 
assign res[86]=in9; 
assign res[87]=in3; 
assign res[88]=neg5; 
assign res[89]=neg10; 
assign res[90]=neg6; 
assign res[91]=neg0; 
assign res[92]=in7; 
assign res[93]=in1; 
assign res[94]=neg3; 
assign res[95]=in12; 
assign res[96]=neg9; 
assign res[97]=neg4; 
assign res[98]=in8; 
assign res[99]=neg12; 
assign res[100]=neg0; 
assign res[101]=neg4; 
assign res[102]=in3; 
assign res[103]=in8; 
assign res[104]=in7; 
assign res[105]=neg7; 
assign res[106]=in7; 
assign res[107]=neg12; 
assign res[108]=neg10; 
assign res[109]=in6; 
assign res[110]=neg4; 
assign res[111]=neg10; 
assign res[112]=neg0; 
assign res[113]=in5; 
assign res[114]=neg7; 
assign res[115]=in12; 
assign res[116]=in3; 
assign res[117]=in8; 
assign res[118]=in12; 
assign res[119]=in7; 
assign res[120]=neg10; 
assign res[121]=in8; 
assign res[122]=neg1; 
assign res[123]=neg6; 
assign res[124]=neg5; 
assign res[125]=in12; 
assign res[126]=in5; 
assign res[127]=in5; 
assign res[128]=neg10; 
assign res[129]=neg13; 
assign res[130]=neg7; 
assign res[131]=in5; 
assign res[132]=neg2; 
assign res[133]=neg7; 
assign res[134]=in9; 
assign res[135]=neg11; 
assign res[136]=neg13; 
assign res[137]=neg13; 
assign res[138]=in6; 
assign res[139]=neg1; 
assign res[140]=neg3; 
assign res[141]=in2; 
assign res[142]=neg13; 
assign res[143]=in12; 
assign res[144]=neg6; 
assign res[145]=in6; 
assign res[146]=neg10; 
assign res[147]=neg4; 
assign res[148]=in2; 
assign res[149]=neg3; 
assign res[150]=in12; 
assign res[151]=in12; 
assign res[152]=neg13; 
assign res[153]=in5; 
assign res[154]=in9; 
assign res[155]=in4; 
assign res[156]=neg1; 
assign res[157]=in2; 
assign res[158]=in6; 
assign res[159]=in1; 
assign res[160]=in11; 
assign res[161]=in5; 
assign res[162]=in7; 
assign res[163]=neg6; 
assign res[164]=neg8; 
assign res[165]=neg7; 
assign res[166]=neg7; 
assign res[167]=neg12; 
assign res[168]=neg3; 
assign res[169]=in12; 
assign res[170]=neg6; 
assign res[171]=neg0; 
assign res[172]=in3; 
assign res[173]=neg13; 
assign res[174]=neg13; 
assign res[175]=in9; 
assign res[176]=in1; 
assign res[177]=neg6; 
assign res[178]=neg1; 
assign res[179]=in12; 
assign res[180]=in1; 
assign res[181]=in6; 
assign res[182]=neg9; 
assign res[183]=in3; 
assign res[184]=neg13; 
assign res[185]=in5; 
assign res[186]=in7; 
assign res[187]=in12; 
assign res[188]=neg5; 
assign res[189]=in9; 
assign res[190]=in3; 
assign res[191]=in11; 
assign res[192]=neg13; 
assign res[193]=in10; 
assign res[194]=neg12; 
assign res[195]=in3; 
assign res[196]=in8; 
assign res[197]=neg6; 
assign res[198]=in6; 
assign res[199]=neg13; 
assign res[200]=neg12; 
assign res[201]=in3; 
assign res[202]=in4; 
assign res[203]=in9; 
assign res[204]=in12; 
assign res[205]=neg6; 
assign res[206]=in12; 
assign res[207]=neg8; 
assign res[208]=neg9; 
assign res[209]=neg4; 
assign res[210]=in3; 
assign res[211]=neg2; 
assign res[212]=in3; 
assign res[213]=neg0; 
assign res[214]=neg3; 
assign res[215]=neg8; 
assign res[216]=in8; 
assign res[217]=in3; 
assign res[218]=neg5; 
assign res[219]=neg4; 
assign res[220]=in11; 
assign res[221]=in10; 
assign res[222]=neg8; 
assign res[223]=in12; 
assign res[224]=in5; 
assign res[225]=neg0; 
assign res[226]=neg1; 
assign res[227]=neg6; 
assign res[228]=neg6; 
assign res[229]=neg11; 
assign res[230]=in12; 
assign res[231]=in7; 
assign res[232]=neg2; 
assign res[233]=in7; 
assign res[234]=neg0; 
assign res[235]=in12; 
assign res[236]=neg8; 
assign res[237]=in2; 
assign res[238]=neg6; 
assign res[239]=in12; 
assign res[240]=neg13; 
assign res[241]=neg8; 
assign res[242]=neg13; 
assign res[243]=neg2; 
assign res[244]=neg8; 
assign res[245]=neg13; 
assign res[246]=neg11; 
assign res[247]=neg0; 
assign res[248]=neg8; 
assign res[249]=neg2; 
assign res[250]=neg4; 
assign res[251]=in1; 
assign res[252]=in1; 
assign res[253]=neg4; 
assign res[254]=neg6; 
assign res[255]=neg11; 
assign res[256]=neg9; 
assign res[257]=in4; 
assign res[258]=in7; 
assign res[259]=in12; 
assign res[260]=in5; 
assign res[261]=in8; 
assign res[262]=neg4; 
assign res[263]=in8; 
assign res[264]=in12; 
assign res[265]=neg13; 
assign res[266]=in7; 
assign res[267]=in12; 
assign res[268]=in2; 
assign res[269]=in7; 
assign res[270]=in11; 
assign res[271]=neg9; 
assign res[272]=in5; 
assign res[273]=neg8; 
assign res[274]=neg4; 
assign res[275]=in9; 
assign res[276]=in9; 
assign res[277]=neg3; 
assign res[278]=neg7; 
assign res[279]=neg12; 
assign res[280]=in5; 
assign res[281]=neg0; 
assign res[282]=in6; 
assign res[283]=in12; 
assign res[284]=in6; 
assign res[285]=neg2; 
assign res[286]=neg10; 
assign res[287]=in10; 
assign res[288]=in1; 
assign res[289]=neg4; 
assign res[290]=neg2; 
assign res[291]=neg13; 
assign res[292]=neg12; 
assign res[293]=in12; 
assign res[294]=neg13; 
assign res[295]=neg6; 
assign res[296]=in1; 
assign res[297]=in3; 
assign res[298]=neg10; 
assign res[299]=neg5; 
assign res[300]=neg13; 
assign res[301]=in1; 
assign res[302]=in5; 
assign res[303]=neg11; 
assign res[304]=neg2; 
assign res[305]=neg7; 
assign res[306]=in9; 
assign res[307]=neg5; 
assign res[308]=in1; 
assign res[309]=in6; 
assign res[310]=neg8; 
assign res[311]=in6; 
assign res[312]=neg4; 
assign res[313]=in1; 
assign res[314]=in11; 
assign res[315]=neg8; 
assign res[316]=in6; 
assign res[317]=neg8; 
assign res[318]=in4; 
assign res[319]=in9; 
assign res[320]=neg5; 
assign res[321]=in3; 
assign res[322]=neg5; 
assign res[323]=in7; 
assign res[324]=neg3; 
assign res[325]=neg8; 
assign res[326]=neg12; 
assign res[327]=in8; 
assign res[328]=neg2; 
assign res[329]=in3; 
assign res[330]=neg13; 
assign res[331]=neg9; 
assign res[332]=neg0; 
assign res[333]=neg5; 
assign res[334]=neg3; 
assign res[335]=in8; 
assign res[336]=neg13; 
assign res[337]=in12; 
assign res[338]=neg8; 
assign res[339]=in9; 
assign res[340]=neg11; 
assign res[341]=neg5; 
assign res[342]=neg2; 
assign res[343]=in11; 
assign res[344]=in9; 
assign res[345]=neg13; 
assign res[346]=neg3; 
assign res[347]=in2; 
assign res[348]=neg13; 
assign res[349]=neg0; 
assign res[350]=in6; 
assign res[351]=neg10; 
assign res[352]=in12; 
assign res[353]=neg7; 
assign res[354]=neg11; 
assign res[355]=in9; 
assign res[356]=neg3; 
assign res[357]=in11; 
assign res[358]=in11; 
assign res[359]=in5; 
assign res[360]=in11; 
assign res[361]=in6; 
assign res[362]=neg5; 
assign res[363]=neg2; 
assign res[364]=in12; 
assign res[365]=in7; 
assign res[366]=neg8; 
assign res[367]=neg2; 
assign res[368]=in1; 
assign res[369]=in7; 
assign res[370]=neg12; 
assign res[371]=neg13; 
assign res[372]=neg2; 
assign res[373]=neg8; 
assign res[374]=in5; 
assign res[375]=neg9; 
assign res[376]=neg1; 
assign res[377]=in5; 
assign res[378]=in7; 
assign res[379]=in10; 
assign res[380]=in5; 
assign res[381]=neg13; 
assign res[382]=neg0; 
assign res[383]=neg13; 
assign res[384]=in12; 
assign res[385]=neg1; 
assign res[386]=neg8; 
assign res[387]=neg9; 
assign res[388]=in11; 
assign res[389]=neg13; 
assign res[390]=neg3; 
assign res[391]=in2; 
assign res[392]=neg10; 
assign res[393]=in12; 
assign res[394]=in1; 
assign res[395]=neg10; 
assign res[396]=neg11; 
assign res[397]=neg6; 
assign res[398]=neg13; 
assign res[399]=neg6; 
assign res[400]=neg13; 
assign res[401]=neg9; 
assign res[402]=neg10; 
assign res[403]=neg7; 
assign res[404]=neg8; 
assign res[405]=neg13; 
assign res[406]=neg6; 
assign res[407]=in5; 
assign res[408]=in12; 
assign res[409]=neg13; 
assign res[410]=in2; 
assign res[411]=neg3; 
assign res[412]=neg13; 
assign res[413]=neg12; 
assign res[414]=neg13; 
assign res[415]=neg1; 
assign res[416]=in9; 
assign res[417]=in3; 
assign res[418]=in3; 
assign res[419]=neg9; 
assign res[420]=in1; 
assign res[421]=in1; 
assign res[422]=in2; 
assign res[423]=neg8; 
assign res[424]=neg10; 
assign res[425]=in9; 
assign res[426]=neg13; 
assign res[427]=in12; 
assign res[428]=neg12; 
assign res[429]=neg5; 
assign res[430]=in2; 
assign res[431]=in7; 
assign res[432]=in6; 
assign res[433]=neg8; 
assign res[434]=in8; 
assign res[435]=neg12; 
assign res[436]=in10; 
assign res[437]=in5; 
assign res[438]=neg9; 
assign res[439]=in9; 
assign res[440]=neg13; 
assign res[441]=in5; 
assign res[442]=neg7; 
assign res[443]=in4; 
assign res[444]=neg2; 
assign res[445]=in3; 
assign res[446]=in2; 
assign res[447]=in12; 
assign res[448]=neg5; 
assign res[449]=in11; 
assign res[450]=neg9; 
assign res[451]=neg13; 
assign res[452]=neg1; 
assign res[453]=in12; 
assign res[454]=neg1; 
assign res[455]=in4; 
assign res[456]=neg0; 
assign res[457]=in6; 
assign res[458]=neg11; 
assign res[459]=in12; 
assign res[460]=neg4; 
assign res[461]=in1; 
assign res[462]=neg6; 
assign res[463]=in1; 
assign res[464]=in7; 
assign res[465]=in1; 
assign res[466]=in12; 
assign res[467]=neg13; 
assign res[468]=neg0; 
assign res[469]=neg13; 
assign res[470]=neg1; 
assign res[471]=in4; 
assign res[472]=in3; 
assign res[473]=neg2; 
assign res[474]=in8; 
assign res[475]=neg3; 
assign res[476]=neg6; 
assign res[477]=neg2; 
assign res[478]=neg9; 
assign res[479]=in10; 
assign res[480]=in7; 
assign res[481]=neg9; 
assign res[482]=neg6; 
assign res[483]=neg1; 
assign res[484]=in5; 
assign res[485]=neg2; 
assign res[486]=neg3; 
assign res[487]=neg8; 
assign res[488]=neg0; 
assign res[489]=in5; 
assign res[490]=in4; 
assign res[491]=in10; 
assign res[492]=neg6; 
assign res[493]=in5; 
assign res[494]=neg0; 
assign res[495]=in5; 
assign res[496]=in8; 
assign res[497]=in11; 
assign res[498]=in9; 
assign res[499]=neg6; 
assign res[500]=neg4; 
assign res[501]=neg12; 
assign res[502]=in4; 
assign res[503]=in9; 
assign res[504]=in3; 
assign res[505]=in4; 
assign res[506]=neg7; 
assign res[507]=neg2; 
assign res[508]=neg0; 
assign res[509]=neg2; 
assign res[510]=neg6; 
assign res[511]=neg11; 
//End Generate ======================================= 

genvar i; 
generate 
for(i=0;i<512;i=i+1) begin : XCon 
	 assign out[i*BW_XCOS +: BW_XCOS] = res[i]; 
end 
endgenerate 

endmodule