module MultX_connect(in0,  in1,  in2,  in3,  in4,  in5,  in6,  in7,  in8, in9, 
		in10, in11, in12, in13, in14, in15, in16, in17, in18, 
		out); 
 
parameter BW_XCOS = 16; 

input signed [BW_XCOS-1:0] in0; 
input signed [BW_XCOS-1:0] in1; 
input signed [BW_XCOS-1:0] in2;  
input signed [BW_XCOS-1:0] in3;  
input signed [BW_XCOS-1:0] in4;  
input signed [BW_XCOS-1:0] in5;  
input signed [BW_XCOS-1:0] in6;  
input signed [BW_XCOS-1:0] in7;  
input signed [BW_XCOS-1:0] in8;  
input signed [BW_XCOS-1:0] in9;  
input signed [BW_XCOS-1:0] in10;  
input signed [BW_XCOS-1:0] in11;  
input signed [BW_XCOS-1:0] in12;  
input signed [BW_XCOS-1:0] in13;  
input signed [BW_XCOS-1:0] in14;  
input signed [BW_XCOS-1:0] in15;
input signed [BW_XCOS-1:0] in16;
input signed [BW_XCOS-1:0] in17;
input signed [BW_XCOS-1:0] in18;

output [512*BW_XCOS-1:0] out; 

wire signed [BW_XCOS-1:0] res [0:511]; 

wire signed [BW_XCOS-1:0] neg0, neg1, neg2, neg3, neg4, neg5,neg6, neg7, neg8, neg9, neg10, neg11, 
	neg12, neg13, neg14, neg15, neg16, neg17, neg18; 

assign neg0=-in0;
assign neg1=-in1; 
assign neg2=-in2; 
assign neg3=-in3; 
assign neg4=-in4; 
assign neg5=-in5; 
assign neg6=-in6; 
assign neg7=-in7; 
assign neg8=-in8; 
assign neg9=-in9; 
assign neg10=-in10; 
assign neg11=-in11; 
assign neg12=-in12; 
assign neg13=-in13; 
assign neg14=-in14; 
assign neg15=-in15; 
assign neg16=-in16;
assign neg17=-in17;
assign neg18=-in18;

//Generating to assign 512 outputs of multiplication == 
assign res[0]=in8; 
assign res[1]=in9; 
assign res[2]=in4; 
assign res[3]=in7; 
assign res[4]=neg11; 
assign res[5]=neg8; 
assign res[6]=in7; 
assign res[7]=in12; 
assign res[8]=in2; 
assign res[9]=in2; 
assign res[10]=in1; 
assign res[11]=in1; 
assign res[12]=neg2; 
assign res[13]=neg2; 
assign res[14]=neg13; 
assign res[15]=neg11; 
assign res[16]=neg13; 
assign res[17]=neg12; 
assign res[18]=in10; 
assign res[19]=in11; 
assign res[20]=neg13; 
assign res[21]=neg8; 
assign res[22]=neg11; 
assign res[23]=neg9; 
assign res[24]=in7; 
assign res[25]=in12; 
assign res[26]=neg4; 
assign res[27]=neg3; 
assign res[28]=neg13; 
assign res[29]=neg12; 
assign res[30]=neg9; 
assign res[31]=neg7; 
assign res[32]=in12; 
assign res[33]=in12; 
assign res[34]=neg3; 
assign res[35]=neg2; 
assign res[36]=neg6; 
assign res[37]=neg4; 
assign res[38]=in11; 
assign res[39]=in12; 
assign res[40]=in4; 
assign res[41]=in5; 
assign res[42]=in5; 
assign res[43]=in10; 
assign res[44]=in3; 
assign res[45]=in6; 
assign res[46]=neg8; 
assign res[47]=neg6; 
assign res[48]=neg2; 
assign res[49]=neg1; 
assign res[50]=neg13; 
assign res[51]=neg8; 
assign res[52]=neg7; 
assign res[53]=neg5; 
assign res[54]=neg4; 
assign res[55]=neg3; 
assign res[56]=neg10; 
assign res[57]=neg6; 
assign res[58]=in5; 
assign res[59]=in6; 
assign res[60]=in5; 
assign res[61]=in7; 
assign res[62]=in1; 
assign res[63]=in4; 
assign res[64]=in9; 
assign res[65]=in11; 
assign res[66]=in4; 
assign res[67]=in4; 
assign res[68]=in2; 
assign res[69]=in4; 
assign res[70]=neg4; 
assign res[71]=neg2; 
assign res[72]=neg8; 
assign res[73]=neg7; 
assign res[74]=in4; 
assign res[75]=in9; 
assign res[76]=neg0; 
assign res[77]=in1; 
assign res[78]=neg13; 
assign res[79]=neg8; 
assign res[80]=neg3; 
assign res[81]=neg2; 
assign res[82]=neg6; 
assign res[83]=neg4; 
assign res[84]=in8; 
assign res[85]=in10; 
assign res[86]=neg0; 
assign res[87]=in1; 
assign res[88]=in7; 
assign res[89]=in11; 
assign res[90]=neg13; 
assign res[91]=neg11; 
assign res[92]=in10; 
assign res[93]=in12; 
assign res[94]=neg6; 
assign res[95]=neg6; 
assign res[96]=in10; 
assign res[97]=in12; 
assign res[98]=neg13; 
assign res[99]=neg8; 
assign res[100]=neg13; 
assign res[101]=neg8; 
assign res[102]=in3; 
assign res[103]=in7; 
assign res[104]=in5; 
assign res[105]=in10; 
assign res[106]=neg1; 
assign res[107]=in1; 
assign res[108]=in3; 
assign res[109]=in5; 
assign res[110]=in2; 
assign res[111]=in3; 
assign res[112]=neg13; 
assign res[113]=neg13; 
assign res[114]=neg13; 
assign res[115]=neg12; 
assign res[116]=neg13; 
assign res[117]=neg11; 
assign res[118]=neg7; 
assign res[119]=neg4; 
assign res[120]=in6; 
assign res[121]=in12; 
assign res[122]=neg9; 
assign res[123]=neg7; 
assign res[124]=neg2; 
assign res[125]=neg0; 
assign res[126]=neg12; 
assign res[127]=neg7; 
assign res[128]=in3; 
assign res[129]=in8; 
assign res[130]=neg7; 
assign res[131]=neg4; 
assign res[132]=neg3; 
assign res[133]=neg1; 
assign res[134]=in2; 
assign res[135]=in5; 
assign res[136]=neg11; 
assign res[137]=neg5; 
assign res[138]=neg1; 
assign res[139]=neg0; 
assign res[140]=in5; 
assign res[141]=in5; 
assign res[142]=neg4; 
assign res[143]=neg4; 
assign res[144]=neg9; 
assign res[145]=neg9; 
assign res[146]=neg12; 
assign res[147]=neg8; 
assign res[148]=in10; 
assign res[149]=in12; 
assign res[150]=in7; 
assign res[151]=in12; 
assign res[152]=neg7; 
assign res[153]=neg6; 
assign res[154]=neg4; 
assign res[155]=neg3; 
assign res[156]=in7; 
assign res[157]=in12; 
assign res[158]=neg7; 
assign res[159]=neg5; 
assign res[160]=neg13; 
assign res[161]=neg12; 
assign res[162]=neg3; 
assign res[163]=neg2; 
assign res[164]=in7; 
assign res[165]=in12; 
assign res[166]=neg13; 
assign res[167]=neg11; 
assign res[168]=in1; 
assign res[169]=in12; 
assign res[170]=in2; 
assign res[171]=in3; 
assign res[172]=neg4; 
assign res[173]=neg2; 
assign res[174]=neg1; 
assign res[175]=in1; 
assign res[176]=in7; 
assign res[177]=in8; 
assign res[178]=in1; 
assign res[179]=in3; 
assign res[180]=in9; 
assign res[181]=in12; 
assign res[182]=neg1; 
assign res[183]=neg1; 
assign res[184]=neg13; 
assign res[185]=neg10; 
assign res[186]=in7; 
assign res[187]=in10; 
assign res[188]=in12; 
assign res[189]=in12; 
assign res[190]=in6; 
assign res[191]=in7; 
assign res[192]=in5; 
assign res[193]=in6; 
assign res[194]=in2; 
assign res[195]=in2; 
assign res[196]=in3; 
assign res[197]=in4; 
assign res[198]=in2; 
assign res[199]=in12; 
assign res[200]=in9; 
assign res[201]=in10; 
assign res[202]=neg8; 
assign res[203]=neg7; 
assign res[204]=neg11; 
assign res[205]=neg4; 
assign res[206]=in1; 
assign res[207]=in2; 
assign res[208]=in6; 
assign res[209]=in7; 
assign res[210]=in2; 
assign res[211]=in3; 
assign res[212]=in6; 
assign res[213]=in11; 
assign res[214]=in3; 
assign res[215]=in8; 
assign res[216]=in7; 
assign res[217]=in9; 
assign res[218]=neg11; 
assign res[219]=neg6; 
assign res[220]=neg10; 
assign res[221]=neg5; 
assign res[222]=neg5; 
assign res[223]=neg3; 
assign res[224]=neg10; 
assign res[225]=neg9; 
assign res[226]=in8; 
assign res[227]=in12; 
assign res[228]=in4; 
assign res[229]=in6; 
assign res[230]=neg10; 
assign res[231]=neg8; 
assign res[232]=in4; 
assign res[233]=in6; 
assign res[234]=neg2; 
assign res[235]=neg2; 
assign res[236]=neg5; 
assign res[237]=neg5; 
assign res[238]=in7; 
assign res[239]=in10; 
assign res[240]=neg9; 
assign res[241]=neg8; 
assign res[242]=neg5; 
assign res[243]=neg5; 
assign res[244]=in8; 
assign res[245]=in9; 
assign res[246]=neg9; 
assign res[247]=neg9; 
assign res[248]=in1; 
assign res[249]=in1; 
assign res[250]=in7; 
assign res[251]=in9; 
assign res[252]=neg2; 
assign res[253]=neg1; 
assign res[254]=in11; 
assign res[255]=in12; 
assign res[256]=neg12; 
assign res[257]=neg6; 
assign res[258]=in3; 
assign res[259]=in7; 
assign res[260]=in5; 
assign res[261]=in10; 
assign res[262]=neg0; 
assign res[263]=in2; 
assign res[264]=neg9; 
assign res[265]=neg5; 
assign res[266]=neg0; 
assign res[267]=in2; 
assign res[268]=neg1; 
assign res[269]=in1; 
assign res[270]=in5; 
assign res[271]=in7; 
assign res[272]=in3; 
assign res[273]=in6; 
assign res[274]=neg13; 
assign res[275]=neg8; 
assign res[276]=neg5; 
assign res[277]=neg3; 
assign res[278]=neg4; 
assign res[279]=neg3; 
assign res[280]=in6; 
assign res[281]=in8; 
assign res[282]=neg7; 
assign res[283]=neg6; 
assign res[284]=neg13; 
assign res[285]=neg5; 
assign res[286]=in1; 
assign res[287]=in3; 
assign res[288]=in4; 
assign res[289]=in8; 
assign res[290]=neg2; 
assign res[291]=in2; 
assign res[292]=in2; 
assign res[293]=in12; 
assign res[294]=neg2; 
assign res[295]=neg0; 
assign res[296]=in4; 
assign res[297]=in9; 
assign res[298]=neg6; 
assign res[299]=neg3; 
assign res[300]=neg3; 
assign res[301]=neg1; 
assign res[302]=in7; 
assign res[303]=in12; 
assign res[304]=in4; 
assign res[305]=in5; 
assign res[306]=neg13; 
assign res[307]=neg9; 
assign res[308]=in7; 
assign res[309]=in8; 
assign res[310]=in7; 
assign res[311]=in7; 
assign res[312]=neg7; 
assign res[313]=neg7; 
assign res[314]=neg8; 
assign res[315]=neg7; 
assign res[316]=neg13; 
assign res[317]=neg12; 
assign res[318]=in2; 
assign res[319]=in3; 
assign res[320]=in10; 
assign res[321]=in12; 
assign res[322]=neg6; 
assign res[323]=neg6; 
assign res[324]=in8; 
assign res[325]=in9; 
assign res[326]=in2; 
assign res[327]=in2; 
assign res[328]=neg11; 
assign res[329]=neg10; 
assign res[330]=neg12; 
assign res[331]=neg7; 
assign res[332]=neg11; 
assign res[333]=neg10; 
assign res[334]=in5; 
assign res[335]=in11; 
assign res[336]=neg2; 
assign res[337]=neg1; 
assign res[338]=neg1; 
assign res[339]=neg0; 
assign res[340]=neg13; 
assign res[341]=neg12; 
assign res[342]=neg10; 
assign res[343]=neg10; 
assign res[344]=neg3; 
assign res[345]=neg2; 
assign res[346]=in2; 
assign res[347]=in3; 
assign res[348]=neg9; 
assign res[349]=neg4; 
assign res[350]=neg4; 
assign res[351]=neg3; 
assign res[352]=neg4; 
assign res[353]=neg2; 
assign res[354]=neg6; 
assign res[355]=neg4; 
assign res[356]=in6; 
assign res[357]=in6; 
assign res[358]=neg13; 
assign res[359]=neg5; 
assign res[360]=in11; 
assign res[361]=in12; 
assign res[362]=in7; 
assign res[363]=in12; 
assign res[364]=neg1; 
assign res[365]=neg0; 
assign res[366]=neg4; 
assign res[367]=neg3; 
assign res[368]=neg7; 
assign res[369]=neg6; 
assign res[370]=neg13; 
assign res[371]=neg8; 
assign res[372]=neg7; 
assign res[373]=neg6; 
assign res[374]=neg8; 
assign res[375]=neg6; 
assign res[376]=neg5; 
assign res[377]=neg4; 
assign res[378]=neg13; 
assign res[379]=neg8; 
assign res[380]=in1; 
assign res[381]=in5; 
assign res[382]=in1; 
assign res[383]=in10; 
assign res[384]=in9; 
assign res[385]=in10; 
assign res[386]=in5; 
assign res[387]=in10; 
assign res[388]=neg1; 
assign res[389]=in1; 
assign res[390]=neg9; 
assign res[391]=neg6; 
assign res[392]=neg1; 
assign res[393]=in1; 
assign res[394]=neg13; 
assign res[395]=neg8; 
assign res[396]=in8; 
assign res[397]=in10; 
assign res[398]=in2; 
assign res[399]=in3; 
assign res[400]=in7; 
assign res[401]=in12; 
assign res[402]=neg10; 
assign res[403]=neg5; 
assign res[404]=neg10; 
assign res[405]=neg8; 
assign res[406]=in4; 
assign res[407]=in8; 
assign res[408]=in3; 
assign res[409]=in8; 
assign res[410]=neg4; 
assign res[411]=neg3; 
assign res[412]=in5; 
assign res[413]=in10; 
assign res[414]=in4; 
assign res[415]=in5; 
assign res[416]=neg9; 
assign res[417]=neg4; 
assign res[418]=neg0; 
assign res[419]=in3; 
assign res[420]=neg12; 
assign res[421]=neg6; 
assign res[422]=in3; 
assign res[423]=in4; 
assign res[424]=neg10; 
assign res[425]=neg10; 
assign res[426]=in8; 
assign res[427]=in12; 
assign res[428]=neg8; 
assign res[429]=neg6; 
assign res[430]=in2; 
assign res[431]=in3; 
assign res[432]=in10; 
assign res[433]=in11; 
assign res[434]=in6; 
assign res[435]=in8; 
assign res[436]=neg7; 
assign res[437]=neg6; 
assign res[438]=neg3; 
assign res[439]=neg3; 
assign res[440]=neg1; 
assign res[441]=neg1; 
assign res[442]=neg3; 
assign res[443]=neg3; 
assign res[444]=neg8; 
assign res[445]=neg8; 
assign res[446]=in4; 
assign res[447]=in12; 
assign res[448]=in2; 
assign res[449]=in3; 
assign res[450]=in6; 
assign res[451]=in11; 
assign res[452]=in3; 
assign res[453]=in7; 
assign res[454]=in11; 
assign res[455]=in12; 
assign res[456]=neg3; 
assign res[457]=neg3; 
assign res[458]=in4; 
assign res[459]=in4; 
assign res[460]=in2; 
assign res[461]=in2; 
assign res[462]=neg10; 
assign res[463]=neg8; 
assign res[464]=neg13; 
assign res[465]=neg11; 
assign res[466]=neg13; 
assign res[467]=neg11; 
assign res[468]=in6; 
assign res[469]=in11; 
assign res[470]=neg0; 
assign res[471]=in1; 
assign res[472]=neg13; 
assign res[473]=neg9; 
assign res[474]=neg9; 
assign res[475]=neg6; 
assign res[476]=neg13; 
assign res[477]=neg8; 
assign res[478]=in5; 
assign res[479]=in8; 
assign res[480]=in2; 
assign res[481]=in3; 
assign res[482]=neg1; 
assign res[483]=neg1; 
assign res[484]=in9; 
assign res[485]=in11; 
assign res[486]=in11; 
assign res[487]=in12; 
assign res[488]=in3; 
assign res[489]=in3; 
assign res[490]=neg1; 
assign res[491]=neg0; 
assign res[492]=in3; 
assign res[493]=in4; 
assign res[494]=neg13; 
assign res[495]=neg10; 
assign res[496]=in5; 
assign res[497]=in12; 
assign res[498]=in8; 
assign res[499]=in9; 
assign res[500]=in7; 
assign res[501]=in8; 
assign res[502]=neg10; 
assign res[503]=neg10; 
assign res[504]=in7; 
assign res[505]=in12; 
assign res[506]=in9; 
assign res[507]=in10; 
assign res[508]=in7; 
assign res[509]=in12; 
assign res[510]=neg1; 
assign res[511]=neg0; 
//End Generate ======================================= 

genvar i; 
generate 
for(i=0;i<512;i=i+1) begin : XCon 
	 assign out[i*BW_XCOS +: BW_XCOS] = res[i]; 
end 
endgenerate 

endmodule
